module lectura_archivo()




endmodule
