`timescale 1ps/1ps;
module tb_FIR_Filter();

initial
 begin
 end
 


endmodule

