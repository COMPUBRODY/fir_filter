
module FIR_Filter(




);


endmodule

