module tb_FIR_Filter();




endmodule

