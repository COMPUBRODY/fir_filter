`timescale 1ps/1ps;

module tb_state_machine()



initial

begin
end

endmodule



