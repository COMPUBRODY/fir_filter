`timescale 1ps/1ps;
module tb_memoria_ram()



initial begin
    
end


endmodule
